`include "defines.sv"

module cpu (
    input logic         Clock,
    input logic         Reset_L,
    input logic         DTAck,
    input logic         IRQ_Timer_H,
    input logic         IRQ_UART_H,
    input logic [31:0]  Instruction,
    input logic [31:0]  DataBus_In,
    output logic        AS_L,
    output logic [3:0]  Byte_Enable,
    output logic        WE_L,
    output logic [31:0] DataBus_Out,
    output logic [31:0] Address,
    output logic        Conduit,
    output logic        Reset_Out
);

    // CPU signals
    enum {LATCH_INSTRUCTION, INITIALIZE, START, WRITE_BACK, INCREMENT_PC, COMPLETE, ACCESS_MEMORY_1, ACCESS_MEMORY_2, WRITE_MEMORY_1, WRITE_MEMORY_2, BRANCH_EQ, BRANCH_NE, BRANCH_LT, BRANCH_GE, BRANCH_LTU, BRANCH_GEU, JUMP_LINK_1, JUMP_LINK_2, JUMP_LINK_3, LOAD_UPPER_IMM_1, CSR_WRITE_BACK, CSRRW_WRITE_1, CSRRW_WRITE_2, CSRRS_WRITE_1, CSRRS_WRITE_2, CSRRC_WRITE_1, CSRRC_WRITE_2, MRET_1, MRET_2, IRQ_1, IRQ_2, IRQ_3, IRQ_4, IRQ_5, CSRRWI_1, CSRRSI_1, CSRRCI_1} State;
    logic           mem_or_reg, jump_link, load_upper_imm, instruction_fetch, save_pc;
    logic           CSR_process;
    logic           CSR_WE_L;
    logic [1:0]     Program_Counter_Increment;
    logic [2:0]     funct3;
    logic [6:0]     funct7, opcode;
    logic [11:0]    imm_I_TYPE, imm_S_TYPE, imm_B_TYPE;
    logic [11:0]    CSR_address;
    logic [19:0]    imm_U_TYPE;
    logic [20:0]    imm_J_TYPE;
    logic [31:0]    datapath_in, Program_Counter, Current_Instruction;
    logic [31:0]    CSR_read_data, CSR_write_data, CSR_read_data_temp;
    logic [31:0]    imm_CSR_TYPE;
    // Data path signals
    logic           reg_bank_write, alu_SRC, negative, overflow, zero;
    logic [3:0]     alu_OP;
    logic [4:0]     rs1, rs2, rd0;
    logic [31:0]    writedata, datapath_out, imm, rs2_output;
    logic MIE, MPIE, MSIE, MTIE, MEIE, MSIP, MTIP, MEIP;
    logic [1:0] MPP, MTVEC_MODE;
    logic [29:0] MTVEC_BASE;
    logic [31:0] MEPC, MCAUSE;

    logic [31:0] MSTATUS_temp;
    logic IRQ_pending;
    logic [31:0]    interrupt_ID;
    logic [11:0]    pending_interrupt_mask;

    datapath HW (
        .clk(Clock),
        .rst_n(Reset_L),
        .write_rb(reg_bank_write),
        .alu_control(alu_OP),
        .alu_source(alu_SRC),
        .rs_1(rs1),
        .rs_2(rs2),
        .rd_0(rd0),
        .writedata(writedata),
        .alu_result(datapath_out),
        .immediate(imm),
        .negative(negative),
        .overflow(overflow),
        .zero(zero),
        .rs2(rs2_output)
    );

    csr CSR (
        .clock(Clock),
        .reset_L(Reset_L),
        .WE_L(CSR_WE_L),
        .address(CSR_address),
        .write_data(CSR_write_data),
        .read_data(CSR_read_data),
        .irq_software(1'b0),
        .irq_timer(IRQ_Timer_H),
        .irq_external(IRQ_UART_H),
        .mstatus_MIE(MIE),
        .mstatus_MPIE(MPIE),
        .mstatus_MPP(MPP),
        .mie_MSIE(MSIE),
        .mie_MTIE(MTIE),
        .mie_MEIE(MEIE),
        .mip_MSIP(MSIP),
        .mip_MTIP(MTIP),
        .mip_MEIP(MEIP),
        .mtvec_MODE(MTVEC_MODE),
        .mtvec_BASE(MTVEC_BASE),
        .mepc_REG(MEPC),
        .mcause_REG(MCAUSE)
    );

    assign datapath_in          = mem_or_reg ? DataBus_In : datapath_out;
    assign rs1                  = Current_Instruction[19:15];
    assign rs2                  = Current_Instruction[24:20];
    assign rd0                  = Current_Instruction[11:7];
    assign funct3               = Current_Instruction[14:12];
    assign funct7               = Current_Instruction[31:25];
    assign opcode               = Current_Instruction[6:0];
    assign imm_I_TYPE           = Current_Instruction[31:20];
    assign imm_S_TYPE           = {Current_Instruction[31:25], Current_Instruction[11:7]}; 
    assign imm_B_TYPE           = {Current_Instruction[31], Current_Instruction[7], Current_Instruction[30:25], Current_Instruction[11:8]};
    assign imm_J_TYPE           = {Current_Instruction[31], Current_Instruction[19:12], Current_Instruction[20], Current_Instruction[30:21], 1'b0};
    assign imm_U_TYPE           = Current_Instruction[31:12];
    assign Address              = instruction_fetch ? Program_Counter : datapath_out;
    //assign CSR_address          = Current_Instruction[31:20];
    assign imm_CSR_TYPE         = {{27{1'b0}}, rs1};
    assign IRQ_pending          = ((MIE == 1'b1) && (((MSIE == 1) && (MSIP == 1)) || ((MTIE == 1) && (MTIP == 1)) || ((MEIE == 1) && (MEIP == 1)))) ? 1'b1 : 1'b0;
    //assign interrupt_ID         = 32'h0;
    assign pending_interrupt_mask   = {MEIP & MEIE, 3'h0, MTIE & MTIP, 3'h0, MSIE & MSIP, 3'h0};

    always @(*) begin
        if (pending_interrupt_mask[11]) begin
            interrupt_ID = 32'd11; // MEIP
        end else if (pending_interrupt_mask[7]) begin
            interrupt_ID = 32'd7; // MTIP
        end else if (pending_interrupt_mask[3]) begin
            interrupt_ID = 32'd3; // MSIP
        end else begin
            interrupt_ID = 32'd0; // no interrupt
        end 
    end
    
    
    always @(*) begin
        case (Byte_Enable) 
            4'b0001: DataBus_Out <= rs2_output;
            4'b0010: DataBus_Out <= rs2_output << 32'd8;
            4'b0100: DataBus_Out <= rs2_output << 32'd16;
            4'b1000: DataBus_Out <= rs2_output << 32'd24;
            4'b0011: DataBus_Out <= rs2_output;
            4'b1100: DataBus_Out <= rs2_output << 32'd16;
            4'b1111: DataBus_Out <= rs2_output;
            default: DataBus_Out <= 32'h00000000;
        endcase
    end
    
    always @(*) begin
        Byte_Enable <= 4'b0000; // disable Byte_Enable by default

        if (funct3 == 3'h0) begin
            case (Address[1:0]) 
                2'b00: Byte_Enable <= 4'b0001; // we are writing a byte at no offset
                2'b01: Byte_Enable <= 4'b0010; // we are writing a byte at offset = 1
                2'b10: Byte_Enable <= 4'b0100; // writing a byte at offset = 2
                2'b11: Byte_Enable <= 4'b1000; // writing a byte at offset = 3
            endcase
        end 

        if (funct3 == 3'h1) begin
            case (Address[1:0]) 
                2'b00: Byte_Enable <= 4'b0011; // writing a half-word at offset = 0
                2'b10: Byte_Enable <= 4'b1100; // writing a half-word at offset = 2
                default: Byte_Enable <= 4'b0000; // we cannot write a half word at offset = 3 or offset = 1, as this is misaligned. Half words must be aligned at byte multiples of 2
            endcase 
        end

        if (funct3 == 3'h2) begin
            Byte_Enable <= 4'b0000; // disable Byte_Enable, unless condition below is met

            if (Address[1:0] == 2'b00) begin
                Byte_Enable <= 4'b1111;
            end
        end
    end

     always @(*) begin
        if (mem_or_reg == 1) begin
            case (funct3)
                3'h0: begin
                    case (Address[1:0])
                        2'b00: writedata <= {{24{datapath_in[7]}}, datapath_in[7:0]};
                        2'b01: writedata <= {{24{datapath_in[15]}}, datapath_in[15:8]};
                        2'b10: writedata <= {{24{datapath_in[23]}}, datapath_in[23:16]};
                        2'b11: writedata <= {{24{datapath_in[31]}}, datapath_in[31:24]};
                    endcase
                end
                3'h1: begin
                    case (Address[1:0])
                        2'b00: writedata <= {{16{datapath_in[15]}}, datapath_in[15:0]};
                        2'b10: writedata <= {{16{datapath_in[31]}}, datapath_in[31:16]};
                        default: writedata <= 32'h00000000;
                    endcase
                end
                3'h2: begin
                    if (Address[1:0] == 2'b00) begin
                        writedata <= datapath_in;
                    end else begin
                        writedata <= 32'h00000000;
                    end
                end
                3'h4: begin
                    case (Address[1:0])
                        2'b00: writedata <= {{24{1'b0}}, datapath_in[7:0]};
                        2'b01: writedata <= {{24{1'b0}}, datapath_in[15:8]};
                        2'b10: writedata <= {{24{1'b0}}, datapath_in[23:16]};
                        2'b11: writedata <= {{24{1'b0}}, datapath_in[31:24]};
                    endcase
                end
                3'h5: begin
                    case (Address[1:0])
                        2'b00: writedata <= {{16{1'b0}}, datapath_in[15:0]};
                        2'b10: writedata <= {{16{1'b0}}, datapath_in[31:16]};
                        default: writedata <= 32'h00000000;
                    endcase
                end
                default: writedata <= 32'h00000000;
            endcase
        end else if (jump_link == 1) begin
            writedata <= Program_Counter + 32'h4;
        end else if (load_upper_imm == 1) begin
            writedata <= imm;
        end else if (CSR_process == 1) begin
            writedata <= CSR_read_data_temp;
        end else begin  
            writedata <= datapath_in;
        end
    end

    always @(posedge Clock, negedge Reset_L) begin
        if (Reset_L == 0) begin
            State                       <= INITIALIZE;
            Program_Counter             <= 32'h00000000;
            AS_L                        <= 1;
            WE_L                        <= 1;
            mem_or_reg                  <= 0;
            alu_OP                      <= 4'h0;
            alu_SRC                     <= 1;
            Conduit                     <= 0;
            jump_link                   <= 0;
            imm                         <= 32'h00000000;
            reg_bank_write              <= 0;
            load_upper_imm              <= 0;
            Conduit                     <= 0;
            Program_Counter_Increment   <= 2'b00;
            Reset_Out                   <= 0;
            instruction_fetch           <= 1;
            CSR_WE_L                    <= 1;
            CSR_process                 <= 0;
            CSR_read_data_temp          <= 32'h0;
            CSR_write_data              <= 32'h0;
            CSR_address                 <= 12'h0;//Current_Instruction[31:20];
            Current_Instruction         <= 32'h00000013; // NOP
        end else begin
            case (State) 
                INITIALIZE: begin
                    State               <= INCREMENT_PC;
                    //Current_Instruction <= Instruction;
                    Reset_Out           <= 1;
                    instruction_fetch   <= 1;
                    save_pc             <= 1;
                end
                START: begin
                    save_pc             <= 0;
                    case (opcode)
                        `R_TYPE: begin
                            State       <= WRITE_BACK;
                            alu_OP      <= {funct7[5], funct3};
                            alu_SRC     <= 1'b1;
                        end
                        `I_TYPE: begin
                            State       <= WRITE_BACK;
                            alu_OP      <= {funct7[5], funct3};
                            alu_SRC     <= 1'b0; 
                            imm         <= {{20{imm_I_TYPE[11]}}, imm_I_TYPE};
                        end       
                        `LOAD_TYPE: begin
                            State       <= ACCESS_MEMORY_1;
                            alu_OP      <= {1'b0, `ADDSUB}; 
                            imm         <= {{20{imm_I_TYPE[11]}}, imm_I_TYPE};
                            alu_SRC     <= 1'b0;
                            instruction_fetch <= 0;
                        end              
                        `S_TYPE: begin
                            State       <= WRITE_MEMORY_1;
                            imm         <= {{20{imm_S_TYPE[11]}}, imm_S_TYPE};
                            alu_SRC     <= 1'b0;
                            alu_OP      <= {1'b0, `ADDSUB};
                            instruction_fetch <= 0;
                        end   
                        `B_TYPE: begin
                            case (funct3)
                                3'h0: begin 
                                        State       <= BRANCH_EQ;
                                        alu_OP      <= {1'b1, `ADDSUB}; 
                                end
                                3'h1: begin
                                        State       <= BRANCH_NE;
                                        alu_OP      <= {1'b1, `ADDSUB};
                                end
                                3'h4: begin 
                                        State       <= BRANCH_LT;
                                        alu_OP      <= {1'b0, `SLT}; // we don't care what the MSB of alu_OP is when using the "set less than" operation    
                                end
                                3'h5: begin 
                                        State       <= BRANCH_GE;
                                        alu_OP      <= {1'b0, `SLT};
                                end
                                3'h6: begin 
                                        State       <= BRANCH_LTU;
                                        alu_OP      <= {1'b0, `SLTU};
                                end
                                3'h7: begin 
                                        State       <= BRANCH_GEU;
                                        alu_OP      <= {1'b0, `SLTU};
                                end
                            endcase
                            alu_SRC     <= 1'b1;
                            imm         <= {{19{imm_B_TYPE[11]}}, imm_B_TYPE, 1'b0};    // zeroth bit of immediate for B-type instructions is always zero (for byte alignment)
                        end
                        `J_TYPE_JAL: begin
                            State           <= JUMP_LINK_1;
                            jump_link       <= 1'b1;
                            imm             <= {{11{imm_J_TYPE[20]}}, imm_J_TYPE};
                        end
                        `J_TYPE_JALR: begin
                            State           <= JUMP_LINK_2;
                            jump_link       <= 1'b1;
                            imm             <= {{20{imm_I_TYPE[11]}}, imm_I_TYPE};
                        end
                        `U_TYPE_LUI: begin
                            State           <= LOAD_UPPER_IMM_1;
                            imm             <= (imm_U_TYPE << 12); 
                            load_upper_imm  <= 1'b1; 
                        end
                        `U_TYPE_AUIPC: begin
                            State           <= LOAD_UPPER_IMM_1;
                            imm             <= (imm_U_TYPE << 12) + Program_Counter;
                            load_upper_imm  <= 1'b1; 
                        end 
                        `CSR_TYPE: begin
                            //CSR_address          <= Current_Instruction[31:20];
                            case (funct3) 
                                `CSRRW: begin
                                    State       <= CSRRW_WRITE_1;
                                    CSR_process <= 1;
                                    CSR_read_data_temp <= CSR_read_data; // save the initial value of whichever CSR we are copying from
                            CSR_address          <= Current_Instruction[31:20];

                                end
                                `CSRRS: begin
                                    State       <= CSRRS_WRITE_1;
                                    CSR_process <= 1;
                                    CSR_read_data_temp <= CSR_read_data;
                            CSR_address          <= Current_Instruction[31:20];

                                end
                                `CSRRC: begin
                                    State       <= CSRRC_WRITE_1;
                                    CSR_process <= 1;
                                    CSR_read_data_temp <= CSR_read_data;
                            CSR_address          <= Current_Instruction[31:20];

                                end
                                `CSRRWI: begin
                                    State       <= CSRRWI_1;
                                    CSR_process <= 1;
                                    // CSR_read_data_temp  <= CSR_read_data;
                                    // CSR_write_data <= imm_CSR_TYPE;
                                    // CSR_WE_L    <= 0;
                            CSR_address          <= Current_Instruction[31:20];

                                end
                                `CSRRSI: begin
                                    State       <= CSRRSI_1;
                                    CSR_process <= 1;
                                    // CSR_read_data_temp  <= CSR_read_data;
                                    // CSR_write_data <= imm_CSR_TYPE | CSR_read_data;
                                    // CSR_WE_L    <= 0;
                            CSR_address          <= Current_Instruction[31:20];

                                end
                                `CSRRCI: begin
                                    State           <= CSRRCI_1;
                                    CSR_process     <= 1;
                                    // CSR_read_data_temp  <= CSR_read_data;
                                    // CSR_write_data  <= CSR_read_data & (~imm_CSR_TYPE);
                                    // CSR_WE_L        <= 0;
                            CSR_address          <= Current_Instruction[31:20];

                                end
                                `MRET: begin
                                    if (Current_Instruction == 32'h30200073) begin
                                        State               <= MRET_1;
                                        CSR_write_data      <= {26'd0, 1'b1, 3'b000, MPIE, 3'b000};
                                        //MSTATUS_temp[3]    <= MPIE;
                                        //MSTATUS_temp[7]     <= 1'b1;
                                        CSR_address <= 12'h300;
                                        //CSR_write_data <= MSTATUS_temp;
                                        CSR_WE_L    <= 1'b1; 
                                    end
                                end
                            endcase
                        end
                        7'b0000000: begin
                            Conduit <= 1'b1;
                            State <= START;
                        end
                        default: State  <= START;
                    endcase
                end
                CSRRCI_1: begin
                    State <= CSR_WRITE_BACK;
                    CSR_read_data_temp  <= CSR_read_data;
                    CSR_write_data  <= CSR_read_data & (~imm_CSR_TYPE);
                    CSR_WE_L        <= 0;
                end
                CSRRSI_1: begin
                    State <= CSR_WRITE_BACK;
                    CSR_read_data_temp  <= CSR_read_data;
                    CSR_write_data <= imm_CSR_TYPE | CSR_read_data;
                    CSR_WE_L    <= 0;
                end
                CSRRWI_1: begin
                    State <= CSR_WRITE_BACK;
                    CSR_read_data_temp  <= CSR_read_data;
                    CSR_write_data <= imm_CSR_TYPE;
                    CSR_WE_L    <= 0;
                end
                MRET_1: begin
                    State <= MRET_2;
                    CSR_WE_L <= 1'b0;

                end
                MRET_2: begin
                    State <= INCREMENT_PC;

                    CSR_WE_L <= 1'b1;
                    Program_Counter <= MEPC;
                end
                CSRRC_WRITE_1: begin
                    State       <= CSRRC_WRITE_2;
                    imm         <= 32'h0;
                    alu_SRC     <= 1'b0;
                    alu_OP      <= {1'b0, `ADDSUB};
                    CSR_read_data_temp <= CSR_read_data;
                end
                CSRRC_WRITE_2: begin
                    State       <= CSR_WRITE_BACK;
                    CSR_write_data <= CSR_read_data_temp & (~datapath_out);
                    CSR_WE_L    <= 0;
                end
                CSRRS_WRITE_1: begin
                    State       <= CSRRS_WRITE_2;
                    imm         <= 32'h0;
                    alu_SRC     <= 1'b0;
                    alu_OP      <= {1'b0, `ADDSUB};
                    CSR_read_data_temp <= CSR_read_data;
                end
                CSRRS_WRITE_2: begin
                    State       <= CSR_WRITE_BACK;
                    CSR_write_data  <= CSR_read_data_temp | datapath_out; 
                    CSR_WE_L    <= 0;
                end
                CSRRW_WRITE_1: begin
                    State       <= CSRRW_WRITE_2;
                    imm         <= 32'h0; // we don't want anything added to whatever is in RS1, ie., RS1 + 0 => output of datapath, to be written back to CSR
                    alu_SRC     <= 1'b0;
                    alu_OP      <= {1'b0, `ADDSUB};
                end
                CSRRW_WRITE_2: begin
                    State       <= CSR_WRITE_BACK;
                    CSR_write_data  <= datapath_out;
                    CSR_WE_L    <= 0;   // write the output of the datapath to CSR
                end
                CSR_WRITE_BACK: begin
                    State       <= COMPLETE;
                    Program_Counter_Increment <= 2'b00;
                    reg_bank_write <= 1;    // writedata bus into datapath and rd0 should be set with CSR data and target destination register, respectively
                    CSR_WE_L    <= 1;
                end
                WRITE_BACK: begin
                    State           <= COMPLETE; 
                    reg_bank_write  <= 1'b1;
                    // increment program counter to next instruction, ie., no jumping
                    //Program_Counter <= Program_Counter + 32'h4;
                    Program_Counter_Increment <= 2'b00;
                end
                COMPLETE: begin
                    if (Program_Counter_Increment == 2'b00) begin
                        // increment program counter by 4
                        Program_Counter <= Program_Counter + 32'h4;
                    end else if (Program_Counter_Increment == 2'b01) begin
                        // increment program counter by immediate
                        Program_Counter <= Program_Counter + imm;
                    end else if (Program_Counter_Increment == 2'b10) begin
                        // set program counter to output of data path
                        Program_Counter <= datapath_out;
                    end

                    if (IRQ_pending == 0) begin
                        State <= INCREMENT_PC;
                        // disable control signals in preparation for next instruction cycle
                        reg_bank_write  <= 1'b0;
                        mem_or_reg      <= 1'b0;
                        WE_L            <= 1'b1;
                        AS_L            <= 1'b1;
                        load_upper_imm  <= 0;
                        instruction_fetch <= 1;
                        jump_link       <= 0;
                        CSR_process     <= 0;
                        // if (Program_Counter_Increment == 2'b00) begin
                        //     // increment program counter by 4
                        //     Program_Counter <= Program_Counter + 32'h4;
                        // end else if (Program_Counter_Increment == 2'b01) begin
                        //     // increment program counter by immediate
                        //     Program_Counter <= Program_Counter + imm;
                        // end else if (Program_Counter_Increment == 2'b10) begin
                        //     // set program counter to output of data path
                        //     Program_Counter <= datapath_out;
                        // end
                    end else begin
                        State               <= IRQ_1;
                        instruction_fetch   <= 1;
                        MSTATUS_temp        <= 32'h0;
                        CSR_write_data      <= Program_Counter;
                        CSR_address         <= 12'h341; 
                        //CSR_WE_L            <= 1'b0;
                    end
                end
                IRQ_1: begin
                    State           <= IRQ_2;
                    //MSTATUS_temp[3] <= 1'b0; // clear MIE bit
                    //MSTATUS_temp[7] <= MIE;     // give MPIE the original value of MIE
                    //CSR_address     <= 12'h300; // mstatus address
                    CSR_WE_L                <= 1'b0; // write to MEPC
                end
                IRQ_2: begin
                    State <= IRQ_3;
                    CSR_write_data      <= {26'd0, MIE, 3'b000, 1'b0, 3'b000};
                    CSR_address         <= 12'h300; // writing to MSTATUS
                    CSR_WE_L            <= 1'b1;
                end
                IRQ_3: begin
                    State <= IRQ_4;
                    //CSR_address         <=12'h342;
                    //CSR_write_data      <= {1'b1, {27{1'b0}}, interrupt_ID[3:0]};
                    CSR_WE_L        <= 1'b0; // write to MSTATUS
                end
                IRQ_4: begin
                    State <= IRQ_5;

                    CSR_address     <= 12'h342; // writing to MCAUSE
                    CSR_write_data  <= {1'b1, 27'b0, interrupt_ID[3:0]};
                    CSR_WE_L    <= 1'b1;
                end
                IRQ_5: begin
                    State <= INCREMENT_PC;
                    CSR_WE_L            <= 1'b0;

                    if (MTVEC_MODE[0] == 1'b0) begin
                        // direct mode 
                        Program_Counter <= {MTVEC_BASE, 2'b00};
                    end else begin
                        // vectored mode 
                        Program_Counter <= {MTVEC_BASE, 2'b00} + (4 * interrupt_ID);
                    end
                end
                INCREMENT_PC: begin
                    State   <= LATCH_INSTRUCTION;
                    // delay one clock cycle for new instruction to appear on output bus of SRAM
                    CSR_WE_L <= 1'b1;
                end
                LATCH_INSTRUCTION: begin
                    State <= START;
                    Current_Instruction <= Instruction;
                    save_pc <= 1;
                end
                ACCESS_MEMORY_1: begin
                    State       <= ACCESS_MEMORY_2;
                    mem_or_reg  <= 1'b1;
                    // WE_L        <= 1'b1;
                    AS_L        <= 1'b0;
                end
                ACCESS_MEMORY_2: begin
                    State           <= DTAck ? COMPLETE : ACCESS_MEMORY_2;
                    reg_bank_write  <= 1'b1;
                    // increment program counter to next instruction, ie., no jumping
                    // Program_Counter <= Program_Counter + 32'h4;
                    Program_Counter_Increment <= 2'b00;
                end
                WRITE_MEMORY_1: begin
                    State       <= WRITE_MEMORY_2;
                    WE_L        <= 1'b0;
                    AS_L        <= 1'b0;
                end
                WRITE_MEMORY_2: begin
                    State <= DTAck ? COMPLETE : WRITE_MEMORY_2;
                    // increment program counter to next instruction, ie., no jumping
                    //Program_Counter <= Program_Counter + 32'h4;
                    Program_Counter_Increment <= 2'b00;
                end
                BRANCH_EQ: begin
                    State   <= COMPLETE;
                    if (zero) begin
                        // add immediate to PC
                        // Program_Counter <= Program_Counter + imm;
                        Program_Counter_Increment <= 2'b01;
                    end else begin
                        // normally increment PC
                        //Program_Counter <= Program_Counter + 32'h4;
                        Program_Counter_Increment <= 2'b00;
                    end
                end
                BRANCH_NE: begin
                    State   <= COMPLETE;
                    if (!zero) begin
                        // increment PC with immediate
                        //Program_Counter <= Program_Counter + imm;
                        Program_Counter_Increment <= 2'b01;
                    end else begin
                        // increment program counter to next instruction
                        //Program_Counter <= Program_Counter + 32'h4;
                        Program_Counter_Increment <= 2'b00;
                    end
                end
                BRANCH_LT: begin
                    State   <= COMPLETE;
                    if (datapath_out == 32'h1) begin // rs1 is less than rs2
                        // increment PC with immediate
                        //Program_Counter <= Program_Counter + imm;
                        Program_Counter_Increment <= 2'b01;
                    end else begin 
                        // increment program counter to next instruction
                        //Program_Counter <= Program_Counter + 32'h4;
                        Program_Counter_Increment <= 2'b00;
                    end 
                end 
                BRANCH_GE: begin
                    State   <= COMPLETE;
                    if (datapath_out == 32'h0) begin
                        // increment PC with immediate
                        //Program_Counter <= Program_Counter + imm;
                        Program_Counter_Increment <= 2'b01;
                    end else begin 
                        // increment program counter to next instruction
                        //Program_Counter <= Program_Counter + 32'h4;
                        Program_Counter_Increment <= 2'b00;
                    end 
                end 
                BRANCH_LTU: begin
                    State   <= COMPLETE;
                    if (datapath_out == 32'h1) begin 
                        // increment PC with immediate
                        //Program_Counter <= Program_Counter + imm;
                        Program_Counter_Increment <= 2'b01;
                    end else begin 
                        // increment program counter to next instruction
                        //Program_Counter <= Program_Counter + 32'h4;
                        Program_Counter_Increment <= 2'b00;
                    end 
                end
                BRANCH_GEU: begin 
                    State   <= COMPLETE;
                    if (datapath_out == 32'h0) begin
                        // increment PC with immediate
                        //Program_Counter <= Program_Counter + imm;
                        Program_Counter_Increment <= 2'b01;
                    end else begin 
                        // increment program counter to next instruction
                        Program_Counter_Increment <= 2'b00;
                        //Program_Counter <= Program_Counter + 32'h4;
                    end 
                end 
                JUMP_LINK_1: begin
                    State           <= COMPLETE;
                    // the writedata line into the datapath (into the register bank) has PC_out + 4 on it, so we just need to set write HIGH
                    reg_bank_write  <= 1'b1; 
                    jump_link       <= 1;
                    // increment program counter with immediate
                    //Program_Counter <= Program_Counter + imm;
                    Program_Counter_Increment <= 2'b01;
                end
                JUMP_LINK_2: begin
                    State           <= JUMP_LINK_3;
                    // write to register bank PC + 4
                    reg_bank_write  <= 1'b1;
                    // disable jump_link so the destination register is not updated after this state
                    jump_link       <= 1'b0;
                    // begin ALU operation to sum RS1 + imm
                    alu_OP[2:0]     <= `ADDSUB;
                    alu_SRC         <= 1'b0;

                end
                JUMP_LINK_3: begin
                    State           <= COMPLETE;

                    // we are no longer writing to the register bank
                    reg_bank_write  <= 0;

                    // program counter gets RS1 + imm
                    //Program_Counter <= datapath_out;
                    Program_Counter_Increment <= 2'b10;
                end
                LOAD_UPPER_IMM_1: begin
                    State           <= COMPLETE; 
                    reg_bank_write  <= 1'b1; // the U-type immediate is on the datapath_in line, just need to write to destination register 
                    // program counter is normally incremented
                    //Program_Counter <= Program_Counter + 32'h4;
                    Program_Counter_Increment <= 2'b00;
                end
            endcase 
        end
    end 
endmodule