module csr (
    input logic         clk,
    input logic         rst_n,
    

);

endmodule: csr