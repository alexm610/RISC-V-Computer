/* opcode */
`define R_TYPE          7'b0110011
`define I_TYPE          7'b0010011
`define S_TYPE          7'b0100011
`define B_TYPE          7'b1100011
`define U_TYPE_LUI      7'b0110111
`define U_TYPE_AUIPC    7'b0010111
`define J_TYPE_JAL      7'b1101111
`define J_TYPE_JALR     7'b1100111
/* ALUop */
`define ADD             4'b0000
`define SUB             4'b0001
`define AND             4'b0010
`define OR              4'b0011
`define NOT             4'b0100 
`define XOR             4'b0101
`define SL              4'b0110
`define SR              4'b0111
