module address_decoder (
        input logic [9:0] address, 
        output logic ROM_Select_H, 
        output logic RAM_Select_H,
        output logic IO_Select_H
);

