// ps2_controller.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module ps2_controller (
		input  wire        address,     //   avalon_ps2_slave.address
		input  wire        chipselect,  //                   .chipselect
		input  wire [3:0]  byteenable,  //                   .byteenable
		input  wire        read,        //                   .read
		input  wire        write,       //                   .write
		input  wire [31:0] writedata,   //                   .writedata
		output wire [31:0] readdata,    //                   .readdata
		output wire        waitrequest, //                   .waitrequest
		input  wire        clk,         //                clk.clk
		inout  wire        PS2_CLK,     // external_interface.CLK
		inout  wire        PS2_DAT,     //                   .DAT
		output wire        irq,         //          interrupt.irq
		input  wire        reset        //              reset.reset
	);

	ps2_controller_ps2_0 ps2_0 (
		.clk         (clk),         //                clk.clk
		.reset       (reset),       //              reset.reset
		.address     (address),     //   avalon_ps2_slave.address
		.chipselect  (chipselect),  //                   .chipselect
		.byteenable  (byteenable),  //                   .byteenable
		.read        (read),        //                   .read
		.write       (write),       //                   .write
		.writedata   (writedata),   //                   .writedata
		.readdata    (readdata),    //                   .readdata
		.waitrequest (waitrequest), //                   .waitrequest
		.irq         (irq),         //          interrupt.irq
		.PS2_CLK     (PS2_CLK),     // external_interface.export
		.PS2_DAT     (PS2_DAT)      //                   .export
	);

endmodule
