/*        ALUop        */
`define ADD 4'b0000
`define SUB 4'b0001
`define AND 4'b0010
`define OR  4'b0011
`define NOT 4'b0100 
`define XOR 4'b0101
`define SL  4'b0110
`define SR  4'b0111
