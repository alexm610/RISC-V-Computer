module memory_1 (input logic clock, input logic reset_n);
    

endmodule: memory_1